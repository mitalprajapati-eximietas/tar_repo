class abc;

	class xyz;

	endclass



endclass
