class seq;




endclass
