










class sequwnce;












endclass
